// Composite Video Timer Verilog Module

// Author: Matthew Knight
// Date: 2017-03-09

// This module takes care of all the timing control for synthesizing a composite
// video signal

module timer();



endmodule
