// Top Module

// Author: Matthew Knight
// Date: 2017-02-22

module spi_comp_top ();

endmodule
